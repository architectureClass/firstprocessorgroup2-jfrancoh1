LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
ENTITY Procesador2_tb IS
END Procesador2_tb;
 
ARCHITECTURE behavior OF Procesador2_tb IS 
 
    COMPONENT Procesador2
    PORT(
         rst : IN  std_logic;
         clk : IN  std_logic;
         cwpc : OUT  std_logic;
         ncwpc : OUT  std_logic;
         nzvcc : OUT  std_logic_vector(3 downto 0);
         resultado : OUT  std_logic_vector(31 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal rst : std_logic := '0';
   signal clk : std_logic := '0';

 	--Outputs
   signal cwpc : std_logic;
   signal ncwpc : std_logic;
   signal nzvcc : std_logic_vector(3 downto 0);
   signal resultado : std_logic_vector(31 downto 0);

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: Procesador2 PORT MAP (
          rst => rst,
          clk => clk,
          cwpc => cwpc,
          ncwpc => ncwpc,
          nzvcc => nzvcc,
          resultado => resultado
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      rst <= '1';
      wait for 100 ns;	
		rst <= '0';
      wait for 100 ns;
      wait for clk_period*10;

      -- insert stimulus here 

      wait;
   end process;

END;
